LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY SUMM IS
GENERIC (N: POSITIVE := 16);
PORT ( IN1: IN SIGNED(N DOWNTO 0);
       IN2: IN SIGNED(N DOWNTO 0);
SUB_ADD: IN STD_LOGIC;
OUTSOM : OUT SIGNED(N DOWNTO 0));
END SUMM;

ARCHITECTURE BEHAV OF SUMM IS
BEGIN
PROCESS (IN1,IN2,SUB_ADD )
BEGIN
IF (SUB_ADD= '0') THEN
OUTSOM<= IN1+IN2;
ELSE
OUTSOM<= IN1-IN2;
END IF;
END PROCESS;
END BEHAV;