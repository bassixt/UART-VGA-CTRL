library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;		 


entity DATAPATH is
port( COM :IN STD_LOGIC_VECTOR(17 DOWNTO 0);
	  ING:IN SIGNED(0 TO 15);
	  CLOCK: IN STD_LOGIC;
      RESET: IN STD_LOGIC;
	  DATA_OUT: OUT SIGNED(15 DOWNTO 0);
	  DONE: OUT STD_LOGIC);
end  DATAPATH ;



architecture behavior of  DATAPATH is

SIGNAL REG_TO_MOL_A,REG_TO_MOL_B,REG_TO_SUM: SIGNED(15 DOWNTO 0);
SIGNAL O_MOL_REG,O_REG_SUM: SIGNED(31 DOWNTO 0);
SIGNAL MUX1_TO_SUM,MUX2_TO_SUM,SUM_TO_REG,REG_TO_REG,REG_TO_MUX2,MUX_TO_MUX:SIGNED(33 DOWNTO 0);


COMPONENT reg_file IS
PORT (  CLOCK: IN STD_LOGIC;
		RESET: IN STD_LOGIC;
		WR_EN: IN STD_LOGIC;
		ADD_A,ADD_B,ADD_C,ADD_IN: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		DATA_A,DATA_B,DATA_C:OUT SIGNED(0 TO 15);
		DATA_IN:IN SIGNED(0 TO 15));
END COMPONENT;


COMPONENT REGN IS
GENERIC (N: POSITIVE := 33);
PORT (R : IN SIGNED(N DOWNTO 0);
	  LOAD: IN STD_LOGIC;
	  ClOCK, RESETN : IN STD_LOGIC;
	  Q : OUT SIGNED(N DOWNTO 0));
END COMPONENT;

COMPONENT SUMM IS
GENERIC (N: POSITIVE := 16);
PORT ( IN1: IN SIGNED(N DOWNTO 0);
       IN2: IN SIGNED(N DOWNTO 0);
SUB_ADD: IN STD_LOGIC;
OUTSOM : OUT SIGNED(N DOWNTO 0));
END COMPONENT;

COMPONENT MUX2TO1 IS
GENERIC( N: POSITIVE :=33);
PORT( I1,I2: IN SIGNED( N DOWNTO 0);
      U: OUT SIGNED (N DOWNTO 0);
      M_SEL: IN STD_LOGIC);
END COMPONENT;


COMPONENT MOLT IS
GENERIC (N: POSITIVE := 15);
PORT ( M1: IN SIGNED(N DOWNTO 0);
       M2: IN SIGNED(N DOWNTO 0);
       SHIFT_MOL: IN STD_LOGIC;
       ClOCK, RESETN ,LDM: IN STD_LOGIC;
       OUTMOL : OUT SIGNED(31 DOWNTO 0));
END COMPONENT;

COMPONENT APPROX IS
PORT (INAPP : IN SIGNED(33 DOWNTO 0);
ClOCK, RESETN ,LD3: IN STD_LOGIC;
OUTAPP: OUT SIGNED(15 DOWNTO 0));
END COMPONENT;
    
BEGIN

RF     :reg_file PORT MAP(CLOCK=>CLOCK,RESET=>RESET,WR_EN=>COM(8),ADD_A=>COM(17 DOWNTO 15),
        ADD_B=>COM(14 DOWNTO 12),ADD_C=>COM(11 DOWNTO 9),ADD_IN=>COM(7 DOWNTO 5),
        DATA_A=>REG_TO_MOL_B,DATA_B=>REG_TO_MOL_A,DATA_C=>REG_TO_SUM,DATA_IN=>ING);                       
REG1  :REGN GENERIC MAP(N=>31)
       PORT MAP( R=>O_MOL_REG,LOAD=>'1',CLOCK=>CLOCK,RESETN=>RESET,Q=>O_REG_SUM);
MOL   :MOLT GENERIC MAP( N=>15)
       PORT MAP ( M1=>REG_TO_MOL_A,M2=>REG_TO_MOL_B,SHIFT_MOL=>COM(4),CLOCK=>CLOCK,RESETN=>RESET,LDM=>'1',OUTMOL=>O_MOL_REG);
SUM   :SUMM GENERIC MAP (N=>33)
       PORT MAP ( IN1=>MUX1_TO_SUM,IN2=>MUX2_TO_SUM,SUB_ADD=>COM(3),OUTSOM=>SUM_TO_REG);
MUX3   : MUX2TO1 GENERIC MAP (N=>33)
       PORT MAP (I2(0)=>'0',I2(1)=>'0',I2(33 DOWNTO 2)=>O_REG_SUM,
       I1(33 DOWNTO 18)=>REG_TO_SUM,I1(17 DOWNTO 0)=>(OTHERS=>'0'),U=>MUX_TO_MUX,M_SEL=>COM(1));
MUX1   : MUX2TO1 GENERIC MAP (N=>33)
       PORT MAP (I2=>MUX_TO_MUX,I1=>REG_TO_MUX2,U=>MUX1_TO_SUM,M_SEL=>COM(2));
MUX2   :MUX2TO1 GENERIC MAP (N=>33)	
        PORT MAP (I1(1)=>'0',I1(0)=>'0',I1(33 DOWNTO 2)=>O_REG_SUM,I2=>REG_TO_MUX2,U=>MUX2_TO_SUM,M_SEL=>COM(1));   
REG2  :REGN GENERIC MAP(N=>33)
       PORT MAP( R=>SUM_TO_REG,LOAD=>'1',CLOCK=>CLOCK,RESETN=>RESET,Q=>REG_TO_REG);
REG3  :REGN GENERIC MAP(N=>33)
       PORT MAP( R=>REG_TO_REG,LOAD=>'1',CLOCK=>CLOCK,RESETN=>RESET,Q=>REG_TO_MUX2);
ROUNDER :APPROX PORT MAP(INAPP=>REG_TO_REG,CLOCK=>CLOCK,RESETN=>RESET,LD3=>'1',OUTAPP=>DATA_OUT);
DONE<=COM(0);
end behavior;