LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY FIFO_CTRL IS
PORT( 	CLOCK,RESETN:IN STD_LOGIC;
		DATA_IN : IN STD_LOGIC_VECTOR(29 DOWNTO 0);
		DATA_OUT: OUT STD_LOGIC_VECTOR(29 DOWNTO 0);
		REQ     : OUT STD_LOGIC;
		POP     : IN STD_LOGIC;
		X       : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
	    Y       : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
		ACK     : IN STD_LOGIC;
		EMPTY   : OUT STD_LOGIC --SEGNALE DI ERRORE
	);
END FIFO_CTRL;

ARCHITECTURE BEHAV OF FIFO_CTRL IS

COMPONENT FIFO IS
GENERIC(CONSTANT N  : positive := 8;  
		CONSTANT M	: positive := 8); 
		
PORT( 	CLOCK,RESETN,PUSH,POP	: IN  STD_LOGIC;
		DATA_IN	   : IN  STD_LOGIC_VECTOR (N-1 DOWNTO 0);
		DATA_OUT   : OUT STD_LOGIC_VECTOR (N-1 DOWNTO 0);
		EMPTY,FULL : OUT STD_LOGIC);
END COMPONENT;

COMPONENT Contatore_Modulo_N IS
GENERIC (N: POSITIVE := 10;
		 M: POSITIVE := 4);
PORT (Data_Input: IN STD_LOGIC_VECTOR(M-1 downto 0);  
	  LD: IN STD_LOGIC;                                    
	  CE: IN STD_LOGIC;
	  INC_DECN: IN STD_LOGIC;							                                     
	  A_RST_n: IN STD_LOGIC;                          
	  CLK: IN STD_LOGIC;                                   
	  Data_Output: BUFFER STD_LOGIC_VECTOR(M-1 downto 0); 
	  TC: OUT STD_LOGIC);   
END COMPONENT;

COMPONENT Contatore_Modulo_N_TC IS
GENERIC (N: POSITIVE := 10;
		 M: POSITIVE := 4);
PORT (Data_Input: IN STD_LOGIC_VECTOR(M-1 downto 0);  
	  LD: IN STD_LOGIC;                                    
	  CE: IN STD_LOGIC; 
	  INC_DECN: IN STD_LOGIC;							                                 
	  A_RST_n: IN STD_LOGIC;                          
	  CLK: IN STD_LOGIC;                                   
	  Data_Output: BUFFER STD_LOGIC_VECTOR(M-1 downto 0); 
	  TC: OUT STD_LOGIC);   
END COMPONENT;

COMPONENT REGN IS
GENERIC (N: POSITIVE := 33);
PORT (R : IN SIGNED(N DOWNTO 0);
LOAD: IN STD_LOGIC;
ClOCK, RESETN : IN STD_LOGIC;
Q : OUT SIGNED(N DOWNTO 0));
END COMPONENT;

TYPE STATE_TYPE IS ( IDLE,START_X,CAMP_W,SAVE_D,TCX_REC,STOP_Y,DEC_1,DEC_2,DEC_3,W_EMPTY);
SIGNAL STATE :STATE_TYPE;
SIGNAL CE_X,CE_Y,CE_PIPE,PUSH,INC_DECN,TCX,FULL:STD_LOGIC;
SIGNAL PI_FI:STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL DATA_OUT_S:STD_LOGIC_VECTOR(7 DOWNTO 0);


BEGIN
TRANSITION: PROCESS( RESETN,CLOCK)
BEGIN
IF RESETN='0' THEN  STATE<= IDLE;
ELSIF ( CLOCK' EVENT AND CLOCK='1') THEN 
CASE STATE IS 
     WHEN IDLE => IF ACK='1' THEN STATE<= START_X; ELSE STATE<= IDLE;END IF;
     WHEN START_X => STATE<= CAMP_W;
     WHEN CAMP_W => STATE<= SAVE_D;
     WHEN SAVE_D => IF FULL='1' THEN STATE<= DEC_1; 
					ELSE 
						IF TCX='1' THEN  STATE<= TCX_REC; 
						ELSE STATE<=SAVE_D; 
						END IF; 
					END IF;
					
     WHEN TCX_REC => STATE<= STOP_Y;
     WHEN STOP_Y => IF FULL='1' THEN STATE<=DEC_1; ELSE STATE<=STOP_Y;END IF;
     WHEN DEC_1=> STATE<=DEC_2;
     WHEN DEC_2=> STATE<=DEC_3;
     WHEN DEC_3=> STATE<=W_EMPTY;
     WHEN W_EMPTY=> IF FULL='0' THEN STATE<= IDLE; ELSE STATE<= W_EMPTY;END IF;
     WHEN OTHERS => STATE <= IDLE;
     END CASE;
 END IF;
 END PROCESS;

 ASM_OUTPUTS: PROCESS( STATE)
BEGIN
REQ<='1';
CE_X<='0';
CE_Y<='0';
CE_PIPE<='1';
INC_DECN<='1';
PUSH<='0';
CASE STATE IS
WHEN IDLE=>
WHEN START_X =>
     CE_X<='1';
WHEN CAMP_W =>
	 CE_X <= '1';
WHEN SAVE_D => 
     CE_X<='1';
     PUSH<='1';  
WHEN TCX_REC => 
     CE_X<='1';
     CE_Y<='1';
     PUSH<='1';
WHEN STOP_Y =>
     CE_X<='1';
     PUSH<='1';
WHEN DEC_1=>
	 CE_X<='1';
	 INC_DECN<='0';
	 REQ<='0';
WHEN DEC_2=>
	 CE_X<='1';
	 INC_DECN<='0';
	 REQ<='0';
WHEN DEC_3=>
	 CE_X<='1';
	 INC_DECN<='0';
	 REQ<='0';	 
WHEN W_EMPTY=>
	 REQ<='0';
END CASE;
END PROCESS;

		--DATA_OUT(7 DOWNTO 6)=>DATA_OUT(21 DOWNTO 20),DATA_OUT(7)=>DATA_OUT(22),DATA_OUT(7)=>DATA_OUT(23)
		--,DATA_OUT(7)=>DATA_OUT(24),DATA_OUT(7)=>DATA_OUT(25),DATA_OUT(7)=>DATA_OUT(26),DATA_OUT(7)=>DATA_OUT(27)
		--,DATA_OUT(7)=>DATA_OUT(28),DATA_OUT(7)=>DATA_OUT(29),DATA_OUT(5 DOWNTO 3)=>DATA_OUT(12 DOWNTO 10)
		--,DATA_OUT(5)=>DATA_OUT(19),DATA_OUT(5)=>DATA_OUT(18),DATA_OUT(5)=>DATA_OUT(17),DATA_OUT(5)=>DATA_OUT(16)
		--,DATA_OUT(5)=>DATA_OUT(15),DATA_OUT(5)=>DATA_OUT(14),DATA_OUT(5)=>DATA_OUT(13),DATA_OUT(2 DOWNTO 0)=>DATA_OUT(2 DOWNTO 0)
		--,DATA_OUT(2)=>DATA_OUT(9),DATA_OUT(2)=>DATA_OUT(8),DATA_OUT(2)=>DATA_OUT(7),DATA_OUT(2)=>DATA_OUT(6),
		--DATA_OUT(2)=>DATA_OUT(5),DATA_OUT(2)=>DATA_OUT(4),DATA_OUT(2)=>DATA_OUT(3)





CONT_TC_638:Contatore_Modulo_N_TC  GENERIC MAP (N=> 640,M=> 10)
       PORT MAP(Data_Input=>"0000000000",LD=>'0',CE=>CE_X,A_RST_n=>RESETN,CLK=>CLOCK,Data_Output=>X,TC=>TCX,INC_DECN=>INC_DECN);      
CONT_480_Y:Contatore_Modulo_N  GENERIC MAP (N=> 480,M=> 9)
       PORT MAP(Data_Input=>"000000000",LD=>'0',CE=>CE_Y,A_RST_n=>RESETN,CLK=>CLOCK,Data_Output=>Y,INC_DECN=>INC_DECN);
PIPE: REGN GENERIC MAP(N=>7)
		PORT MAP (R=>SIGNED(DATA_IN(7 DOWNTO 0)),LOAD=>CE_PIPE,CLOCK=>CLOCK,RESETN=>RESETN,STD_LOGIC_VECTOR(Q)=>PI_FI);
FIFO_MEM: FIFO GENERIC MAP(N=>8,M=>16)
		PORT MAP (CLOCK=>CLOCK,RESETN=>RESETN,PUSH=>PUSH,POP=>POP,DATA_IN=>PI_FI,
		DATA_OUT=>DATA_OUT_S,EMPTY=>EMPTY,FULL=>FULL);
DATA_OUT(7 DOWNTO 0)<=DATA_OUT_S;
DATA_OUT(8)<=DATA_OUT_S(7);
DATA_OUT(9)<=DATA_OUT_S(7);
DATA_OUT(10)<=DATA_OUT_S(7);
DATA_OUT(11)<=DATA_OUT_S(7);
DATA_OUT(12)<=DATA_OUT_S(7);
DATA_OUT(13)<=DATA_OUT_S(7);
DATA_OUT(14)<=DATA_OUT_S(7);
DATA_OUT(15)<=DATA_OUT_S(7);
DATA_OUT(16)<=DATA_OUT_S(7);
DATA_OUT(17)<=DATA_OUT_S(7);
DATA_OUT(18)<=DATA_OUT_S(7);
DATA_OUT(19)<=DATA_OUT_S(7);
DATA_OUT(20)<=DATA_OUT_S(7);
DATA_OUT(21)<=DATA_OUT_S(7);
DATA_OUT(22)<=DATA_OUT_S(7);
DATA_OUT(23)<=DATA_OUT_S(7);
DATA_OUT(24)<=DATA_OUT_S(7);
DATA_OUT(25)<=DATA_OUT_S(7);
DATA_OUT(26)<=DATA_OUT_S(7);
DATA_OUT(27)<=DATA_OUT_S(7);
DATA_OUT(28)<=DATA_OUT_S(7);
DATA_OUT(29)<=DATA_OUT_S(7);		
END BEHAV;