LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY STATUS_PLA IS
PORT ( 
CC,STATUS,LSB_IN : IN STD_LOGIC;
LSB_OUT : OUT STD_LOGIC);
END STATUS_PLA;
ARCHITECTURE Behavior OF STATUS_PLA IS
BEGIN
LSB_OUT<=( CC AND STATUS) OR ( NOT CC AND LSB_IN);
END Behavior;