LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY APPROX IS

PORT (INAPP : IN SIGNED(33 DOWNTO 0);
ClOCK, RESETN ,LD3: IN STD_LOGIC;
OUTAPP: OUT SIGNED(15 DOWNTO 0));
END APPROX;

ARCHITECTURE BEHAV OF APPROX IS

COMPONENT REGN IS
GENERIC (N: POSITIVE := 33);
PORT (R : IN SIGNED(N DOWNTO 0);
LOAD: IN STD_LOGIC;
ClOCK, RESETN : IN STD_LOGIC;
Q : OUT SIGNED(N DOWNTO 0));
END COMPONENT;

COMPONENT MUX2TO1 IS
GENERIC( N: POSITIVE :=33);
PORT( I1,I2: IN SIGNED( N DOWNTO 0);
      U: OUT SIGNED (N DOWNTO 0);
      M_SEL: IN STD_LOGIC);
END COMPONENT;

COMPONENT SUMM IS
GENERIC (N: POSITIVE := 16);
PORT ( IN1: IN SIGNED(N DOWNTO 0);
       IN2: IN SIGNED(N DOWNTO 0);
SUB_ADD: IN STD_LOGIC;
OUTSOM : OUT SIGNED(N DOWNTO 0));
END COMPONENT;

SIGNAL OUTAND: STD_LOGIC ;
SIGNAL OUTMUX1: SIGNED(16 DOWNTO 0);
SIGNAL OUTS: SIGNED(16 DOWNTO 0);

BEGIN



OUTAND<=INAPP(17) AND NOT INAPP(16) AND NOT INAPP(15) AND NOT INAPP(14) AND NOT INAPP(13) AND NOT INAPP(12) AND NOT INAPP(11)
        AND NOT INAPP(10) AND NOT INAPP(9) AND NOT INAPP(8) AND NOT INAPP(7) AND NOT INAPP(6) AND NOT INAPP(5) AND NOT INAPP(4)
        AND NOT INAPP(3) AND NOT INAPP(2) AND NOT INAPP(1) AND NOT INAPP(0);

SUM1:SUMM GENERIC MAP (N=>16)
     PORT MAP(IN1=>INAPP(33 DOWNTO 17), IN2=>"00000000000000001", SUB_ADD=>'0',OUTSOM=>OUTS);
     
MUX1: MUX2TO1 GENERIC MAP (N=>16)
      PORT MAP(I1=>OUTS, I2(16 DOWNTO 2)=>OUTS(16 DOWNTO 2),I2(1)=>'0',I2(0)=>OUTS(0),M_SEL=>OUTAND,U=>OUTMUX1);   

REG16:REGN GENERIC MAP (N=>15)
       PORT MAP(R=>OUTMUX1(16 DOWNTO 1),LOAD=>LD3,RESETN=>RESETN,CLOCK=>CLOCK,Q=>OUTAPP);
END BEHAV;