library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;		 


entity VGASINCR is
port( 
	   CLK,RESETN,EMPTY: IN STD_LOGIC;
	   VGA_CLOCK,VGA_SINK,VGA_BLANK,VGA_VS,VGA_HS,POP : OUT STD_LOGIC );
end  VGASINCR ;

ARCHITECTURE BEHAV OF VGASINCR IS


COMPONENT Cont797 IS
PORT (                                   
	  CE1: IN STD_LOGIC;                                  
	  RESETN: IN STD_LOGIC;                             
	  CLK: IN STD_LOGIC;                                   
	  OUTCON: OUT UNSIGNED(9 downto 0); 
	  TC94: OUT STD_LOGIC;
	  TC141: OUT STD_LOGIC;
	  TC781: OUT STD_LOGIC;
	  TC796: OUT STD_LOGIC);                                  
END COMPONENT;

COMPONENT Cont524 IS
PORT (                                   
	  CE2: IN STD_LOGIC;                                  
	  RESETN: IN STD_LOGIC;                             
	  CLK: IN STD_LOGIC;                                   
	  OUTCON2: OUT UNSIGNED(9 downto 0); 
	  TCL1: OUT STD_LOGIC;
	  TCL34: OUT STD_LOGIC;
	  TCL514: OUT STD_LOGIC;
	  TCL524: OUT STD_LOGIC);                                  
END CoMPONENT;

TYPE STATE_TYPE IS ( IDLE,CE1_VA,CE2_VA,CE1_VB,CE2_VB,CE1_HA,CE1_HB,AUS_1,CE1_HC,AUS_2,CE1_HD,CE2_VC,CE1_VD,CE2_VD);
TYPE STATE_TYPE2 IS ( IDLE2,CE1_HA2,CE1_HB2,AUS_12,CE1_HC2,AUS_22,CE2_VC2,CE1_HD2);

SIGNAL STATE :STATE_TYPE;
SIGNAL STATE2 :STATE_TYPE2;

SIGNAL CE1,CE2,TC94,TC141,TC781,TC796,TCL1,TCL34,TCL514,TCL524: STD_LOGIC;
SIGNAL OUTCON1:UNSIGNED(9 downto 0); 
SIGNAL OUTCON2: UNSIGNED(9 downto 0); 
BEGIN 
TRANSITION_VERTICAL: PROCESS( RESETN, CLK)
BEGIN
IF RESETN='0' THEN  STATE<= IDLE;
ELSIF ( CLK' EVENT AND CLK='1') THEN 
CASE STATE IS 
     WHEN IDLE => IF EMPTY='1' THEN STATE<=IDLE; ELSE STATE<=CE1_VA;END IF;
     WHEN CE1_VA => IF TC796='1' THEN STATE<=CE2_VA ; ELSE STATE<= CE1_VA;END IF;
     WHEN CE2_VA => IF TCL1='1' THEN STATE<=CE1_VB ; ELSE STATE<= CE1_VA;END IF;
     WHEN CE1_VB => IF TC796='1' THEN STATE<=CE2_VB ; ELSE STATE<= CE1_VB;END IF;
     WHEN CE2_VB => IF TCL34='1' THEN STATE<=CE1_HA ; ELSE STATE<= CE1_VB;END IF;
     WHEN CE1_HA => IF TC94='1' THEN STATE<=CE1_HB ; ELSE STATE<= CE1_HA;END IF;
     WHEN CE1_HB=> IF TC141='1' THEN STATE<=AUS_1; ELSE STATE<= CE1_HB;END IF;
     WHEN AUS_1=> STATE<=CE1_HC;
     WHEN CE1_HC => IF TC781='1' THEN STATE<=AUS_2; ELSE STATE<= CE1_HC;END IF;
     WHEN AUS_2=> STATE<=CE1_HD;
     WHEN CE1_HD => IF TC796='1' THEN STATE<=CE2_VC ; ELSE STATE<= CE1_HD;END IF;
     WHEN CE2_VC => IF TCL514='1' THEN STATE<=CE1_VD ; ELSE STATE<= CE1_HA;END IF;
     WHEN CE1_VD => IF TC796='1' THEN STATE<=CE2_VD ; ELSE STATE<= CE1_VD;END IF;
     WHEN CE2_VD => IF TCL524='1' THEN STATE<=CE1_VA; ELSE STATE<= CE1_VD;END IF;
     
     END CASE;
    END IF;
 END PROCESS;
 
ASM_OUTPUTS_VERTICAL: PROCESS( STATE)
BEGIN

CE2<='0';
VGA_SINK<='0';
VGA_BLANK<='0';
VGA_VS<='1';

POP<='0';

CASE STATE IS
WHEN IDLE=>
WHEN CE1_VA =>
 
     VGA_VS<='0';
WHEN CE2_VA=>
 
     CE2<='1';
     VGA_VS<='0';
WHEN CE1_VB =>   

WHEN CE2_VB =>

     CE2<='1';
WHEN CE1_HA =>

WHEN CE1_HB=> 
  
WHEN AUS_1=> 
   
     POP<='1';
WHEN CE1_HC=>
   
     VGA_BLANK<='1';
   
     POP<='1';
WHEN AUS_2=>

     VGA_BLANK<='1';

WHEN CE1_HD =>

WHEN CE2_VC=>

     CE2<='1';
WHEN CE1_VD =>

WHEN CE2_VD =>

     CE2<='1';
  
      END CASE;
 END PROCESS;
 -------------------------
 
 
 
 TRANSITION_HOR: PROCESS( RESETN, CLK)
BEGIN
IF RESETN='0' THEN  STATE2<= IDLE2;
ELSIF ( CLK' EVENT AND CLK='1') THEN 
CASE STATE2 IS 
     WHEN IDLE2 => IF EMPTY='1' THEN STATE2<=IDLE2; ELSE STATE2<=CE1_HA2;END IF;
     WHEN CE1_HA2 => IF TC94='1' THEN STATE2<=CE1_HB2 ; ELSE STATE2<= CE1_HA2;END IF;
     WHEN CE1_HB2=> IF TC141='1' THEN STATE2<=AUS_12; ELSE STATE2<= CE1_HB2;END IF;
     WHEN AUS_12=> STATE2<=CE1_HC2;
     WHEN CE1_HC2 => IF TC781='1' THEN STATE2<=AUS_22; ELSE STATE2<= CE1_HC2;END IF;
     WHEN AUS_22=> STATE2<=CE1_HD2;
     WHEN CE1_HD2 => IF TC796='1' THEN STATE2<=CE2_VC2 ; ELSE STATE2<= CE1_HD2;END IF;
     WHEN CE2_VC2 => STATE2<=CE1_HA2;
     WHEN OTHERS=> STATE2<=IDLE2;
    END CASE;
    END IF;
 END PROCESS;
 
ASM_OUTPUTS_HOR: PROCESS( STATE2)
BEGIN
CE1<='0';

VGA_HS<='1';


CASE STATE2 IS
WHEN IDLE2=>
WHEN CE1_HA2 =>
     CE1<='1';
     VGA_HS<='0';
WHEN CE1_HB2=> 
     CE1<='1';
WHEN AUS_12=> 
     CE1<='1';
  
WHEN CE1_HC2=>
     CE1<='1';
   
WHEN AUS_22=>
     CE1<='1';
  
WHEN CE1_HD2 =>
     CE1<='1';
WHEN CE2_VC2=>
     CE1<='1';

      END CASE;
 END PROCESS;
 
 VGA_CLOCK<=CLK;
 
 CONTATORE797: Cont797 port map ( CE1=>CE1, RESETN=>RESETN,CLK=>CLK,OUTCON=>OUTCON1,TC94=>TC94,TC141=>TC141,TC781=>TC781,TC796=>TC796);
 CONTATORE524: Cont524 port map ( CE2=>CE2, RESETN=>RESETN,CLK=>CLK,OUTCON2=>OUTCON2,TCL1=>TCL1,TCL34=>TCL34,TCL514=>TCL514,TCL524=>TCL524); 
     
     
END BEHAV;
     
     