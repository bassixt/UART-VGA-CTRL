library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;		 


entity butterfly is
port( DATA_IN: IN SIGNED(15 DOWNTO 0);
	  START,CLK,RESETN : IN STD_LOGIC;
	  DATA_OUT: OUT SIGNED(15 DOWNTO 0);
	  DONE : OUT STD_LOGIC
	 );
end  butterfly ;

architecture behavior of  butterfly is

SIGNAL ADDR_UROM: STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL ROM_TO_UIR: STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL UIR_OUT: STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL PLA_TO_SEQ: STD_LOGIC;


COMPONENT microrom is
port(	
		ADDR	: in std_logic_vector(4 downto 0);
		DATA_OUT: out STD_LOGIC_VECTOR(23 downto 0));
END COMPONENT;

COMPONENT REGN_STD IS
GENERIC (N: POSITIVE := 33);
PORT (R : IN STD_LOGIC_VECTOR(N DOWNTO 0);
LOAD: IN STD_LOGIC;
ClOCK, RESETN : IN STD_LOGIC;
Q : OUT STD_LOGIC_VECTOR(N DOWNTO 0));
END COMPONENT;

COMPONENT STATUS_PLA IS
PORT ( 
CC,STATUS,LSB_IN : IN STD_LOGIC;
LSB_OUT : OUT STD_LOGIC);
END COMPONENT;

COMPONENT REGN_F_STD IS
GENERIC (N: POSITIVE := 33);
PORT (R : IN STD_LOGIC_VECTOR(N DOWNTO 0);
LOAD: IN STD_LOGIC;
ClOCK, RESETN : IN STD_LOGIC;
Q : OUT STD_LOGIC_VECTOR(N DOWNTO 0));
END COMPONENT;

COMPONENT DATAPATH is
port( COM :IN STD_LOGIC_VECTOR(17 DOWNTO 0);
	  ING:IN SIGNED(0 TO 15);
	  CLOCK: IN STD_LOGIC;
      RESET: IN STD_LOGIC;
	  DATA_OUT: OUT SIGNED(15 DOWNTO 0);
	  DONE: OUT STD_LOGIC);
end  COMPONENT ;




    
BEGIN

MUROM:microrom PORT MAP(ADDR=>ADDR_UROM,DATA_OUT=>ROM_TO_UIR);

MUIR   :REGN_F_STD GENERIC MAP(N=>23)  
		     PORT MAP(R=>ROM_TO_UIR,LOAD=>'1',ClOCK=>CLK, RESETN=>RESETN,Q=>UIR_OUT);
		     
MUPC   :REGN_STD GENERIC MAP(N=>4)
		     PORT MAP(R(4 DOWNTO 1)=>UIR_OUT(22 DOWNTO 19),R(0)=>PLA_TO_SEQ,LOAD=>'1',ClOCK=>CLK, RESETN=>RESETN,Q=>ADDR_UROM);
		     
S_PLA  :STATUS_PLA  PORT MAP (CC=>UIR_OUT(23),STATUS=>START,LSB_IN=>UIR_OUT(18),LSB_OUT=>PLA_TO_SEQ);

DP     : DATAPATH PORT MAP(COM=>UIR_OUT(17 DOWNTO 0),ING=>DATA_IN,CLOCK=>CLK,RESET=>RESETN,DATA_OUT=>DATA_OUT,DONE=>DONE);

end behavior;

