LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY MUX2TO1 IS
GENERIC( N: POSITIVE :=33);
PORT(I1,I2: IN SIGNED( N DOWNTO 0);
     U: OUT SIGNED (N DOWNTO 0);
     M_SEL: IN STD_LOGIC);
END MUX2TO1;

ARCHITECTURE BEHAV OF MUX2TO1 IS
BEGIN 
MUXPROCESS: PROCESS(I1,I2,M_SEL)
BEGIN
IF M_SEL = '0' THEN
	U <= I1;
ELSE
	U <= I2;
END IF;
END PROCESS;
END BEHAV;