LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY reg_file IS
PORT (  CLOCK: IN STD_LOGIC;
		RESET: IN STD_LOGIC;
		WR_EN: IN STD_LOGIC;
		ADD_A,ADD_B,ADD_C,ADD_IN: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		DATA_A,DATA_B,DATA_C:OUT SIGNED(0 TO 15);
		DATA_IN:IN SIGNED(0 TO 15));
END reg_file;

ARCHITECTURE BEHAVIOR OF reg_file IS

TYPE REG IS ARRAY (0 TO 4) OF SIGNED(15 DOWNTO 0);
SIGNAL DATA: REG;
BEGIN 
MEM: PROCESS(RESET,CLOCK)
BEGIN
IF RESET = '0' THEN
		DATA<=(OTHERS => "0000000000000000");
ELSIF CLOCK' EVENT AND CLOCK='1' THEN
	  IF WR_EN = '1'THEN
		DATA(to_integer(unsigned(ADD_IN)))<=DATA_IN;

	  END IF;
END IF;
END PROCESS;

DATA_A<=DATA(to_integer(unsigned(ADD_A)));
DATA_B<=DATA(to_integer(unsigned(ADD_B)));
DATA_C<=DATA(to_integer(unsigned(ADD_C)));
END ARCHITECTURE;